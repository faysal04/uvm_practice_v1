package mux_pkg;
  import uvm_pkg::*;
  `include "uvm_macros.svh"

  //`include "mux_intf.sv";
  `include "mux_tx.sv";
  `include "mux_seq.sv";
  `include "mux_sequencer.sv";
  `include "mux_driver.sv";
  `include "mux_monitor.sv";
  `include "mux_agent.sv";
  `include "mux_env.sv";
  `include "mux_test.sv";

endpackage : mux_pkg