class mux_seq extends uvm_sequence#(mux_tx);

  `uvm_object_utils(mux_seq)

  mux_tx txn;

  function new (string name="mux_seq");
    super.new(name);
  endfunction

  virtual task body();
    txn=mux_tx::type_id::create("txn");
    repeat(100) begin
      start_item(txn);
      txn.randomizee;
      finish_item(txn);
    end
  endtask

endclass
