package mux_pkg;
  `include "mux_intf.sv";
  `include "mux_tx.sv";
  `include "mux_seq.sv";
  `include "mux_sequencer.sv";
  `include "mux_driver.sv";
  `include "mux_moitor.sv";
  `include "mux_agent.sv";
  `include "mux_env.sv";
  `include "mux_test.sv";
  `include "top.sv";
endpackage : mux_pkg